magic
tech sky130A
magscale 1 2
timestamp 1729243200
<< nwell >>
rect -178 -106 822 2824
<< nsubdiff >>
rect -142 2754 -82 2788
rect 726 2754 786 2788
rect -142 2728 -108 2754
rect 752 2728 786 2754
rect -142 -36 -108 -10
rect 752 -36 786 -10
rect -142 -70 -82 -36
rect 726 -70 786 -36
<< nsubdiffcont >>
rect -82 2754 726 2788
rect -142 -10 -108 2728
rect 752 -10 786 2728
rect -82 -70 726 -36
<< poly >>
rect -58 2716 34 2732
rect -58 2682 -42 2716
rect -8 2682 34 2716
rect -58 2666 34 2682
rect 4 2634 34 2666
rect 608 2690 700 2706
rect 608 2656 650 2690
rect 684 2656 700 2690
rect 608 2640 700 2656
rect 608 2634 638 2640
rect -58 2008 34 2024
rect -58 1974 -42 2008
rect -8 1974 34 2008
rect 92 1996 292 2112
rect -58 1958 34 1974
rect 4 1900 34 1958
rect 608 1984 700 2000
rect 608 1950 650 1984
rect 684 1950 700 1984
rect 608 1934 700 1950
rect 608 1900 638 1934
rect 94 1286 550 1404
rect 6 738 36 796
rect -56 722 36 738
rect -56 688 -40 722
rect -6 688 36 722
rect 610 758 640 790
rect 610 742 702 758
rect 610 708 652 742
rect 686 708 702 742
rect -56 672 36 688
rect 352 580 552 696
rect 610 692 702 708
rect 6 52 36 84
rect -56 37 36 52
rect -56 3 -40 37
rect -6 3 36 37
rect -56 -14 36 3
rect 610 52 640 84
rect 610 36 702 52
rect 610 2 652 36
rect 686 2 702 36
rect 610 -14 702 2
<< polycont >>
rect -42 2682 -8 2716
rect 650 2656 684 2690
rect -42 1974 -8 2008
rect 650 1950 684 1984
rect -40 688 -6 722
rect 652 708 686 742
rect -40 3 -6 37
rect 652 2 686 36
<< locali >>
rect -142 2754 -82 2788
rect 726 2754 786 2788
rect -142 2728 -108 2754
rect 752 2728 786 2754
rect -58 2682 -42 2716
rect -8 2682 8 2716
rect -42 2608 -8 2682
rect 634 2656 650 2690
rect 684 2656 700 2690
rect 650 2608 684 2656
rect -58 1974 -42 2008
rect -8 1974 8 2008
rect -42 1900 -8 1974
rect 634 1950 650 1984
rect 684 1950 700 1984
rect 650 1900 684 1950
rect -40 722 -6 796
rect 652 742 686 790
rect -56 688 -40 722
rect -6 688 10 722
rect 636 708 652 742
rect 686 708 702 742
rect -40 37 -6 84
rect 652 36 686 84
rect -56 2 -40 36
rect -6 2 10 36
rect 636 2 652 36
rect 686 2 702 36
rect -142 -36 -108 -10
rect 752 -36 786 -10
rect -142 -70 -82 -36
rect 726 -70 786 -36
<< viali >>
rect 650 2754 684 2788
rect -42 2682 -8 2716
rect 650 2656 684 2690
rect -42 1974 -8 2008
rect 650 1950 684 1984
rect -40 688 -6 722
rect 652 708 686 742
rect -40 3 -6 36
rect -40 2 -6 3
rect 652 2 686 36
rect -40 -70 -6 -36
<< metal1 >>
rect 638 2788 696 2794
rect 638 2754 650 2788
rect 684 2754 696 2788
rect -54 2716 4 2722
rect -54 2682 -42 2716
rect -8 2682 4 2716
rect -54 2676 4 2682
rect 638 2690 696 2754
rect -48 2608 -2 2676
rect 638 2656 650 2690
rect 684 2656 696 2690
rect 638 2650 696 2656
rect 644 2608 690 2650
rect -48 2596 88 2608
rect -62 2220 -52 2596
rect 0 2220 88 2596
rect -48 2208 88 2220
rect 300 2166 344 2608
rect 556 2208 692 2608
rect 556 2166 600 2208
rect 300 2122 600 2166
rect -54 2008 4 2014
rect -54 1974 -42 2008
rect -8 1974 4 2008
rect -54 1968 4 1974
rect -48 1900 -2 1968
rect -46 1888 90 1900
rect -46 1512 36 1888
rect 88 1512 98 1888
rect -46 1500 90 1512
rect 122 1410 262 1462
rect 44 1228 264 1280
rect 44 1192 86 1228
rect -46 792 90 1192
rect -46 728 0 792
rect -52 722 6 728
rect -52 688 -40 722
rect -6 688 6 722
rect -52 682 6 688
rect 300 570 344 2122
rect 638 1984 696 1990
rect 638 1950 650 1984
rect 684 1950 696 1984
rect 638 1944 696 1950
rect 644 1894 690 1944
rect 556 1506 692 1894
rect 380 1458 520 1462
rect 556 1458 602 1506
rect 380 1414 602 1458
rect 380 1410 520 1414
rect 382 1228 522 1280
rect 554 1178 690 1180
rect 544 802 554 1178
rect 606 802 690 1178
rect 554 792 690 802
rect 646 748 692 790
rect 640 742 698 748
rect 640 708 652 742
rect 686 708 698 742
rect 640 702 698 708
rect 42 526 344 570
rect 42 484 86 526
rect -46 84 90 484
rect 300 84 344 526
rect 558 96 642 472
rect 694 96 704 472
rect 558 84 694 96
rect -46 42 0 84
rect 646 42 692 84
rect -52 36 6 42
rect -52 2 -40 36
rect -6 2 6 36
rect -52 -36 6 2
rect 640 36 698 42
rect 640 2 652 36
rect 686 2 698 36
rect 640 -4 698 2
rect -52 -70 -40 -36
rect -6 -70 6 -36
rect -52 -76 6 -70
<< via1 >>
rect -52 2220 0 2596
rect 36 1512 88 1888
rect 554 802 606 1178
rect 642 96 694 472
<< metal2 >>
rect -52 2596 0 2606
rect -52 2095 0 2220
rect -56 2086 0 2095
rect 638 2088 698 2097
rect -56 2021 0 2030
rect 627 2028 636 2088
rect 698 2028 705 2088
rect -52 664 0 2021
rect 638 2019 698 2028
rect 36 1888 88 1898
rect 36 1372 88 1512
rect 36 1318 606 1372
rect 554 1178 606 1318
rect 554 792 606 802
rect 639 664 697 2019
rect -65 604 -56 664
rect 4 604 13 664
rect 638 662 698 664
rect 638 606 640 662
rect 696 606 698 662
rect 638 472 698 606
rect 638 450 642 472
rect 694 450 698 472
rect 642 86 694 96
<< via2 >>
rect -56 2030 0 2086
rect 636 2028 698 2088
rect -56 604 4 664
rect 640 606 696 662
<< metal3 >>
rect -61 2088 5 2091
rect 631 2088 703 2093
rect -61 2086 636 2088
rect -61 2030 -56 2086
rect 0 2030 636 2086
rect -61 2028 636 2030
rect 698 2028 703 2088
rect -61 2025 5 2028
rect 631 2023 703 2028
rect -61 664 9 669
rect 635 664 701 667
rect -61 604 -56 664
rect 4 662 701 664
rect 4 606 640 662
rect 696 606 701 662
rect 4 604 701 606
rect -61 599 9 604
rect 635 601 701 604
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729224599
transform 1 0 623 0 1 2408
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729224599
transform 1 0 623 0 1 1700
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729224599
transform 1 0 625 0 1 990
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729224599
transform 1 0 19 0 1 2408
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729224599
transform 1 0 19 0 1 1700
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729224599
transform 1 0 625 0 1 284
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729224599
transform 1 0 21 0 1 990
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729224599
transform 1 0 21 0 1 284
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729223976
transform 1 0 321 0 1 2408
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729223976
transform 1 0 321 0 1 1700
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729223976
transform 1 0 323 0 1 990
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729223976
transform 1 0 323 0 1 284
box -323 -300 323 300
<< labels >>
flabel metal1 668 2726 668 2726 0 FreeSans 800 0 0 0 VDD
port 4 nsew
flabel space 58 1400 58 1400 0 FreeSans 800 0 0 0 D1
port 5 nsew
flabel metal1 574 1440 574 1440 0 FreeSans 800 0 0 0 D2
port 6 nsew
flabel space 666 1340 666 1340 0 FreeSans 800 0 0 0 D5
port 7 nsew
<< end >>
